// main.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module main (
		input  wire       arbitro_0_conduit_end_beginbursttransfer,   //            arbitro_0_conduit_end.beginbursttransfer
		output wire       arbitro_0_conduit_end_writeresponsevalid_n, //                                 .writeresponsevalid_n
		input  wire       button_down_external_connection_export,     //  button_down_external_connection.export
		output wire       button_enter_external_connection_export,    // button_enter_external_connection.export
		input  wire       button_exit_external_connection_export,     //  button_exit_external_connection.export
		input  wire       button_up_external_connection_export,       //    button_up_external_connection.export
		input  wire       clk_clk,                                    //                              clk.clk
		output wire       lcd_output_external_RS,                     //              lcd_output_external.RS
		output wire       lcd_output_external_RW,                     //                                 .RW
		inout  wire [7:0] lcd_output_external_data,                   //                                 .data
		output wire       lcd_output_external_E,                      //                                 .E
		output wire       led_b_external_connection_export,           //        led_b_external_connection.export
		output wire       led_g_external_connection_export,           //        led_g_external_connection.export
		output wire       led_r_external_connection_export,           //        led_r_external_connection.export
		input  wire       uart_main_external_connection_rxd,          //    uart_main_external_connection.rxd
		output wire       uart_main_external_connection_txd           //                                 .txd
	);

	wire         nios2_processor_jtag_debug_module_reset_reset;                                     // nios2_processor:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller:reset_in1]
	wire         nios2_processor_custom_instruction_master_readra;                                  // nios2_processor:D_ci_readra -> nios2_processor_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] nios2_processor_custom_instruction_master_a;                                       // nios2_processor:D_ci_a -> nios2_processor_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] nios2_processor_custom_instruction_master_b;                                       // nios2_processor:D_ci_b -> nios2_processor_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] nios2_processor_custom_instruction_master_c;                                       // nios2_processor:D_ci_c -> nios2_processor_custom_instruction_master_translator:ci_slave_c
	wire         nios2_processor_custom_instruction_master_readrb;                                  // nios2_processor:D_ci_readrb -> nios2_processor_custom_instruction_master_translator:ci_slave_readrb
	wire  [31:0] nios2_processor_custom_instruction_master_ipending;                                // nios2_processor:W_ci_ipending -> nios2_processor_custom_instruction_master_translator:ci_slave_ipending
	wire   [7:0] nios2_processor_custom_instruction_master_n;                                       // nios2_processor:D_ci_n -> nios2_processor_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] nios2_processor_custom_instruction_master_result;                                  // nios2_processor_custom_instruction_master_translator:ci_slave_result -> nios2_processor:E_ci_result
	wire         nios2_processor_custom_instruction_master_estatus;                                 // nios2_processor:W_ci_estatus -> nios2_processor_custom_instruction_master_translator:ci_slave_estatus
	wire  [31:0] nios2_processor_custom_instruction_master_datab;                                   // nios2_processor:E_ci_datab -> nios2_processor_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] nios2_processor_custom_instruction_master_dataa;                                   // nios2_processor:E_ci_dataa -> nios2_processor_custom_instruction_master_translator:ci_slave_dataa
	wire         nios2_processor_custom_instruction_master_writerc;                                 // nios2_processor:D_ci_writerc -> nios2_processor_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] nios2_processor_custom_instruction_master_translator_comb_ci_master_result;        // nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_result -> nios2_processor_custom_instruction_master_translator:comb_ci_master_result
	wire         nios2_processor_custom_instruction_master_translator_comb_ci_master_readra;        // nios2_processor_custom_instruction_master_translator:comb_ci_master_readra -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] nios2_processor_custom_instruction_master_translator_comb_ci_master_a;             // nios2_processor_custom_instruction_master_translator:comb_ci_master_a -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] nios2_processor_custom_instruction_master_translator_comb_ci_master_b;             // nios2_processor_custom_instruction_master_translator:comb_ci_master_b -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         nios2_processor_custom_instruction_master_translator_comb_ci_master_readrb;        // nios2_processor_custom_instruction_master_translator:comb_ci_master_readrb -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] nios2_processor_custom_instruction_master_translator_comb_ci_master_c;             // nios2_processor_custom_instruction_master_translator:comb_ci_master_c -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         nios2_processor_custom_instruction_master_translator_comb_ci_master_estatus;       // nios2_processor_custom_instruction_master_translator:comb_ci_master_estatus -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] nios2_processor_custom_instruction_master_translator_comb_ci_master_ipending;      // nios2_processor_custom_instruction_master_translator:comb_ci_master_ipending -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] nios2_processor_custom_instruction_master_translator_comb_ci_master_datab;         // nios2_processor_custom_instruction_master_translator:comb_ci_master_datab -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] nios2_processor_custom_instruction_master_translator_comb_ci_master_dataa;         // nios2_processor_custom_instruction_master_translator:comb_ci_master_dataa -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         nios2_processor_custom_instruction_master_translator_comb_ci_master_writerc;       // nios2_processor_custom_instruction_master_translator:comb_ci_master_writerc -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] nios2_processor_custom_instruction_master_translator_comb_ci_master_n;             // nios2_processor_custom_instruction_master_translator:comb_ci_master_n -> nios2_processor_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_result;         // nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_result -> nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_readra;         // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_readra -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_a;              // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_a -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_b;              // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_b -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_readrb;         // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_readrb -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_c;              // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_c -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_estatus;        // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_estatus -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_ipending;       // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_ipending -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_datab;          // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_datab -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_dataa;          // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_dataa -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_writerc;        // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_writerc -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_n;              // nios2_processor_custom_instruction_master_comb_xconnect:ci_master0_n -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] nios2_processor_custom_instruction_master_comb_slave_translator0_ci_master_result; // arbitro_0:result -> nios2_processor_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] nios2_processor_custom_instruction_master_comb_slave_translator0_ci_master_datab;  // nios2_processor_custom_instruction_master_comb_slave_translator0:ci_master_datab -> arbitro_0:datab
	wire  [31:0] nios2_processor_custom_instruction_master_comb_slave_translator0_ci_master_dataa;  // nios2_processor_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> arbitro_0:dataa
	wire  [31:0] nios2_processor_data_master_readdata;                                              // mm_interconnect_0:nios2_processor_data_master_readdata -> nios2_processor:d_readdata
	wire         nios2_processor_data_master_waitrequest;                                           // mm_interconnect_0:nios2_processor_data_master_waitrequest -> nios2_processor:d_waitrequest
	wire         nios2_processor_data_master_debugaccess;                                           // nios2_processor:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_processor_data_master_debugaccess
	wire  [15:0] nios2_processor_data_master_address;                                               // nios2_processor:d_address -> mm_interconnect_0:nios2_processor_data_master_address
	wire   [3:0] nios2_processor_data_master_byteenable;                                            // nios2_processor:d_byteenable -> mm_interconnect_0:nios2_processor_data_master_byteenable
	wire         nios2_processor_data_master_read;                                                  // nios2_processor:d_read -> mm_interconnect_0:nios2_processor_data_master_read
	wire         nios2_processor_data_master_write;                                                 // nios2_processor:d_write -> mm_interconnect_0:nios2_processor_data_master_write
	wire  [31:0] nios2_processor_data_master_writedata;                                             // nios2_processor:d_writedata -> mm_interconnect_0:nios2_processor_data_master_writedata
	wire  [31:0] nios2_processor_instruction_master_readdata;                                       // mm_interconnect_0:nios2_processor_instruction_master_readdata -> nios2_processor:i_readdata
	wire         nios2_processor_instruction_master_waitrequest;                                    // mm_interconnect_0:nios2_processor_instruction_master_waitrequest -> nios2_processor:i_waitrequest
	wire  [15:0] nios2_processor_instruction_master_address;                                        // nios2_processor:i_address -> mm_interconnect_0:nios2_processor_instruction_master_address
	wire         nios2_processor_instruction_master_read;                                           // nios2_processor:i_read -> mm_interconnect_0:nios2_processor_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                          // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                       // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                              // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                             // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire   [7:0] mm_interconnect_0_lcd_output_control_slave_readdata;                               // lcd_output:readdata -> mm_interconnect_0:lcd_output_control_slave_readdata
	wire   [1:0] mm_interconnect_0_lcd_output_control_slave_address;                                // mm_interconnect_0:lcd_output_control_slave_address -> lcd_output:address
	wire         mm_interconnect_0_lcd_output_control_slave_read;                                   // mm_interconnect_0:lcd_output_control_slave_read -> lcd_output:read
	wire         mm_interconnect_0_lcd_output_control_slave_begintransfer;                          // mm_interconnect_0:lcd_output_control_slave_begintransfer -> lcd_output:begintransfer
	wire         mm_interconnect_0_lcd_output_control_slave_write;                                  // mm_interconnect_0:lcd_output_control_slave_write -> lcd_output:write
	wire   [7:0] mm_interconnect_0_lcd_output_control_slave_writedata;                              // mm_interconnect_0:lcd_output_control_slave_writedata -> lcd_output:writedata
	wire  [31:0] mm_interconnect_0_nios2_processor_jtag_debug_module_readdata;                      // nios2_processor:jtag_debug_module_readdata -> mm_interconnect_0:nios2_processor_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest;                   // nios2_processor:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_processor_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess;                   // mm_interconnect_0:nios2_processor_jtag_debug_module_debugaccess -> nios2_processor:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_processor_jtag_debug_module_address;                       // mm_interconnect_0:nios2_processor_jtag_debug_module_address -> nios2_processor:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_read;                          // mm_interconnect_0:nios2_processor_jtag_debug_module_read -> nios2_processor:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable;                    // mm_interconnect_0:nios2_processor_jtag_debug_module_byteenable -> nios2_processor:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_processor_jtag_debug_module_write;                         // mm_interconnect_0:nios2_processor_jtag_debug_module_write -> nios2_processor:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_processor_jtag_debug_module_writedata;                     // mm_interconnect_0:nios2_processor_jtag_debug_module_writedata -> nios2_processor:jtag_debug_module_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                                  // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                                    // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                     // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                                  // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                                       // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                                   // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                                       // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_led_r_s1_chipselect;                                             // mm_interconnect_0:led_r_s1_chipselect -> led_r:chipselect
	wire  [31:0] mm_interconnect_0_led_r_s1_readdata;                                               // led_r:readdata -> mm_interconnect_0:led_r_s1_readdata
	wire   [1:0] mm_interconnect_0_led_r_s1_address;                                                // mm_interconnect_0:led_r_s1_address -> led_r:address
	wire         mm_interconnect_0_led_r_s1_write;                                                  // mm_interconnect_0:led_r_s1_write -> led_r:write_n
	wire  [31:0] mm_interconnect_0_led_r_s1_writedata;                                              // mm_interconnect_0:led_r_s1_writedata -> led_r:writedata
	wire  [31:0] mm_interconnect_0_button_exit_s1_readdata;                                         // button_exit:readdata -> mm_interconnect_0:button_exit_s1_readdata
	wire   [1:0] mm_interconnect_0_button_exit_s1_address;                                          // mm_interconnect_0:button_exit_s1_address -> button_exit:address
	wire         mm_interconnect_0_button_enter_s1_chipselect;                                      // mm_interconnect_0:button_enter_s1_chipselect -> button_enter:chipselect
	wire  [31:0] mm_interconnect_0_button_enter_s1_readdata;                                        // button_enter:readdata -> mm_interconnect_0:button_enter_s1_readdata
	wire   [1:0] mm_interconnect_0_button_enter_s1_address;                                         // mm_interconnect_0:button_enter_s1_address -> button_enter:address
	wire         mm_interconnect_0_button_enter_s1_write;                                           // mm_interconnect_0:button_enter_s1_write -> button_enter:write_n
	wire  [31:0] mm_interconnect_0_button_enter_s1_writedata;                                       // mm_interconnect_0:button_enter_s1_writedata -> button_enter:writedata
	wire  [31:0] mm_interconnect_0_button_down_s1_readdata;                                         // button_down:readdata -> mm_interconnect_0:button_down_s1_readdata
	wire   [1:0] mm_interconnect_0_button_down_s1_address;                                          // mm_interconnect_0:button_down_s1_address -> button_down:address
	wire         mm_interconnect_0_led_b_s1_chipselect;                                             // mm_interconnect_0:led_b_s1_chipselect -> led_b:chipselect
	wire  [31:0] mm_interconnect_0_led_b_s1_readdata;                                               // led_b:readdata -> mm_interconnect_0:led_b_s1_readdata
	wire   [1:0] mm_interconnect_0_led_b_s1_address;                                                // mm_interconnect_0:led_b_s1_address -> led_b:address
	wire         mm_interconnect_0_led_b_s1_write;                                                  // mm_interconnect_0:led_b_s1_write -> led_b:write_n
	wire  [31:0] mm_interconnect_0_led_b_s1_writedata;                                              // mm_interconnect_0:led_b_s1_writedata -> led_b:writedata
	wire         mm_interconnect_0_led_g_s1_chipselect;                                             // mm_interconnect_0:led_g_s1_chipselect -> led_g:chipselect
	wire  [31:0] mm_interconnect_0_led_g_s1_readdata;                                               // led_g:readdata -> mm_interconnect_0:led_g_s1_readdata
	wire   [1:0] mm_interconnect_0_led_g_s1_address;                                                // mm_interconnect_0:led_g_s1_address -> led_g:address
	wire         mm_interconnect_0_led_g_s1_write;                                                  // mm_interconnect_0:led_g_s1_write -> led_g:write_n
	wire  [31:0] mm_interconnect_0_led_g_s1_writedata;                                              // mm_interconnect_0:led_g_s1_writedata -> led_g:writedata
	wire         mm_interconnect_0_uart_main_s1_chipselect;                                         // mm_interconnect_0:uart_main_s1_chipselect -> uart_main:chipselect
	wire  [15:0] mm_interconnect_0_uart_main_s1_readdata;                                           // uart_main:readdata -> mm_interconnect_0:uart_main_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_main_s1_address;                                            // mm_interconnect_0:uart_main_s1_address -> uart_main:address
	wire         mm_interconnect_0_uart_main_s1_read;                                               // mm_interconnect_0:uart_main_s1_read -> uart_main:read_n
	wire         mm_interconnect_0_uart_main_s1_begintransfer;                                      // mm_interconnect_0:uart_main_s1_begintransfer -> uart_main:begintransfer
	wire         mm_interconnect_0_uart_main_s1_write;                                              // mm_interconnect_0:uart_main_s1_write -> uart_main:write_n
	wire  [15:0] mm_interconnect_0_uart_main_s1_writedata;                                          // mm_interconnect_0:uart_main_s1_writedata -> uart_main:writedata
	wire  [31:0] mm_interconnect_0_button_up_s1_readdata;                                           // button_up:readdata -> mm_interconnect_0:button_up_s1_readdata
	wire   [1:0] mm_interconnect_0_button_up_s1_address;                                            // mm_interconnect_0:button_up_s1_address -> button_up:address
	wire         irq_mapper_receiver0_irq;                                                          // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                          // uart_main:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_processor_d_irq_irq;                                                         // irq_mapper:sender_irq -> nios2_processor:d_irq
	wire         rst_controller_reset_out_reset;                                                    // rst_controller:reset_out -> [arbitro_0:reset, button_down:reset_n, button_enter:reset_n, button_exit:reset_n, button_up:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, lcd_output:reset_n, led_b:reset_n, led_g:reset_n, led_r:reset_n, mm_interconnect_0:nios2_processor_reset_n_reset_bridge_in_reset_reset, nios2_processor:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, uart_main:reset_n]
	wire         rst_controller_reset_out_reset_req;                                                // rst_controller:reset_req -> [nios2_processor:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	arbitro arbitro_0 (
		.clk    (clk_clk),                                                                           //                         clock.clk
		.reset  (rst_controller_reset_out_reset),                                                    //                         reset.reset
		.start  (),                                                                                  // nios_custom_instruction_slave.start
		.dataa  (nios2_processor_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  //                              .dataa
		.datab  (nios2_processor_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //                              .datab
		.result (nios2_processor_custom_instruction_master_comb_slave_translator0_ci_master_result), //                              .result
		.done   (),                                                                                  //                              .done
		.rx     (arbitro_0_conduit_end_beginbursttransfer),                                          //                   conduit_end.beginbursttransfer
		.tx     (arbitro_0_conduit_end_writeresponsevalid_n)                                         //                              .writeresponsevalid_n
	);

	main_button_down button_down (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_button_down_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_down_s1_readdata), //                    .readdata
		.in_port  (button_down_external_connection_export)     // external_connection.export
	);

	main_button_enter button_enter (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_button_enter_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_enter_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_enter_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_enter_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_enter_s1_readdata),   //                    .readdata
		.out_port   (button_enter_external_connection_export)       // external_connection.export
	);

	main_button_down button_exit (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_button_exit_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_exit_s1_readdata), //                    .readdata
		.in_port  (button_exit_external_connection_export)     // external_connection.export
	);

	main_button_down button_up (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address  (mm_interconnect_0_button_up_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_up_s1_readdata), //                    .readdata
		.in_port  (button_up_external_connection_export)     // external_connection.export
	);

	main_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	main_lcd_output lcd_output (
		.reset_n       (~rst_controller_reset_out_reset),                          //         reset.reset_n
		.clk           (clk_clk),                                                  //           clk.clk
		.begintransfer (mm_interconnect_0_lcd_output_control_slave_begintransfer), // control_slave.begintransfer
		.read          (mm_interconnect_0_lcd_output_control_slave_read),          //              .read
		.write         (mm_interconnect_0_lcd_output_control_slave_write),         //              .write
		.readdata      (mm_interconnect_0_lcd_output_control_slave_readdata),      //              .readdata
		.writedata     (mm_interconnect_0_lcd_output_control_slave_writedata),     //              .writedata
		.address       (mm_interconnect_0_lcd_output_control_slave_address),       //              .address
		.LCD_RS        (lcd_output_external_RS),                                   //      external.export
		.LCD_RW        (lcd_output_external_RW),                                   //              .export
		.LCD_data      (lcd_output_external_data),                                 //              .export
		.LCD_E         (lcd_output_external_E)                                     //              .export
	);

	main_button_enter led_b (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_led_b_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_b_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_b_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_b_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_b_s1_readdata),   //                    .readdata
		.out_port   (led_b_external_connection_export)       // external_connection.export
	);

	main_button_enter led_g (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_led_g_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_g_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_g_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_g_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_g_s1_readdata),   //                    .readdata
		.out_port   (led_g_external_connection_export)       // external_connection.export
	);

	main_button_enter led_r (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_led_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_r_s1_readdata),   //                    .readdata
		.out_port   (led_r_external_connection_export)       // external_connection.export
	);

	main_nios2_processor nios2_processor (
		.clk                                   (clk_clk),                                                         //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                              //                          .reset_req
		.d_address                             (nios2_processor_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_processor_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_processor_data_master_read),                                //                          .read
		.d_readdata                            (nios2_processor_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_processor_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_processor_data_master_write),                               //                          .write
		.d_writedata                           (nios2_processor_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_processor_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_processor_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_processor_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_processor_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_processor_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_processor_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_processor_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_processor_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_processor_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_processor_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_processor_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_processor_jtag_debug_module_writedata),   //                          .writedata
		.E_ci_result                           (nios2_processor_custom_instruction_master_result),                // custom_instruction_master.result
		.D_ci_a                                (nios2_processor_custom_instruction_master_a),                     //                          .a
		.D_ci_b                                (nios2_processor_custom_instruction_master_b),                     //                          .b
		.D_ci_c                                (nios2_processor_custom_instruction_master_c),                     //                          .c
		.D_ci_n                                (nios2_processor_custom_instruction_master_n),                     //                          .n
		.D_ci_readra                           (nios2_processor_custom_instruction_master_readra),                //                          .readra
		.D_ci_readrb                           (nios2_processor_custom_instruction_master_readrb),                //                          .readrb
		.D_ci_writerc                          (nios2_processor_custom_instruction_master_writerc),               //                          .writerc
		.E_ci_dataa                            (nios2_processor_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_datab                            (nios2_processor_custom_instruction_master_datab),                 //                          .datab
		.E_ci_multi_clock                      (),                                                                //                          .clk
		.E_ci_multi_reset                      (),                                                                //                          .reset
		.E_ci_multi_reset_req                  (),                                                                //                          .reset_req
		.W_ci_estatus                          (nios2_processor_custom_instruction_master_estatus),               //                          .estatus
		.W_ci_ipending                         (nios2_processor_custom_instruction_master_ipending)               //                          .ipending
	);

	main_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	main_uart_main uart_main (
		.clk           (clk_clk),                                      //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address       (mm_interconnect_0_uart_main_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_main_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_main_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_main_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_main_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_main_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_main_s1_readdata),      //                    .readdata
		.rxd           (uart_main_external_connection_rxd),            // external_connection.export
		.txd           (uart_main_external_connection_txd),            //                    .export
		.irq           (irq_mapper_receiver1_irq)                      //                 irq.irq
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) nios2_processor_custom_instruction_master_translator (
		.ci_slave_dataa            (nios2_processor_custom_instruction_master_dataa),                              //       ci_slave.dataa
		.ci_slave_datab            (nios2_processor_custom_instruction_master_datab),                              //               .datab
		.ci_slave_result           (nios2_processor_custom_instruction_master_result),                             //               .result
		.ci_slave_n                (nios2_processor_custom_instruction_master_n),                                  //               .n
		.ci_slave_readra           (nios2_processor_custom_instruction_master_readra),                             //               .readra
		.ci_slave_readrb           (nios2_processor_custom_instruction_master_readrb),                             //               .readrb
		.ci_slave_writerc          (nios2_processor_custom_instruction_master_writerc),                            //               .writerc
		.ci_slave_a                (nios2_processor_custom_instruction_master_a),                                  //               .a
		.ci_slave_b                (nios2_processor_custom_instruction_master_b),                                  //               .b
		.ci_slave_c                (nios2_processor_custom_instruction_master_c),                                  //               .c
		.ci_slave_ipending         (nios2_processor_custom_instruction_master_ipending),                           //               .ipending
		.ci_slave_estatus          (nios2_processor_custom_instruction_master_estatus),                            //               .estatus
		.comb_ci_master_dataa      (nios2_processor_custom_instruction_master_translator_comb_ci_master_dataa),    // comb_ci_master.dataa
		.comb_ci_master_datab      (nios2_processor_custom_instruction_master_translator_comb_ci_master_datab),    //               .datab
		.comb_ci_master_result     (nios2_processor_custom_instruction_master_translator_comb_ci_master_result),   //               .result
		.comb_ci_master_n          (nios2_processor_custom_instruction_master_translator_comb_ci_master_n),        //               .n
		.comb_ci_master_readra     (nios2_processor_custom_instruction_master_translator_comb_ci_master_readra),   //               .readra
		.comb_ci_master_readrb     (nios2_processor_custom_instruction_master_translator_comb_ci_master_readrb),   //               .readrb
		.comb_ci_master_writerc    (nios2_processor_custom_instruction_master_translator_comb_ci_master_writerc),  //               .writerc
		.comb_ci_master_a          (nios2_processor_custom_instruction_master_translator_comb_ci_master_a),        //               .a
		.comb_ci_master_b          (nios2_processor_custom_instruction_master_translator_comb_ci_master_b),        //               .b
		.comb_ci_master_c          (nios2_processor_custom_instruction_master_translator_comb_ci_master_c),        //               .c
		.comb_ci_master_ipending   (nios2_processor_custom_instruction_master_translator_comb_ci_master_ipending), //               .ipending
		.comb_ci_master_estatus    (nios2_processor_custom_instruction_master_translator_comb_ci_master_estatus),  //               .estatus
		.ci_slave_multi_clk        (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_reset      (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_clken      (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_reset_req  (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_start      (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_done       (),                                                                             //    (terminated)
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                         //    (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                         //    (terminated)
		.ci_slave_multi_result     (),                                                                             //    (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                                  //    (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                         //    (terminated)
		.ci_slave_multi_a          (5'b00000),                                                                     //    (terminated)
		.ci_slave_multi_b          (5'b00000),                                                                     //    (terminated)
		.ci_slave_multi_c          (5'b00000),                                                                     //    (terminated)
		.multi_ci_master_clk       (),                                                                             //    (terminated)
		.multi_ci_master_reset     (),                                                                             //    (terminated)
		.multi_ci_master_clken     (),                                                                             //    (terminated)
		.multi_ci_master_reset_req (),                                                                             //    (terminated)
		.multi_ci_master_start     (),                                                                             //    (terminated)
		.multi_ci_master_done      (1'b0),                                                                         //    (terminated)
		.multi_ci_master_dataa     (),                                                                             //    (terminated)
		.multi_ci_master_datab     (),                                                                             //    (terminated)
		.multi_ci_master_result    (32'b00000000000000000000000000000000),                                         //    (terminated)
		.multi_ci_master_n         (),                                                                             //    (terminated)
		.multi_ci_master_readra    (),                                                                             //    (terminated)
		.multi_ci_master_readrb    (),                                                                             //    (terminated)
		.multi_ci_master_writerc   (),                                                                             //    (terminated)
		.multi_ci_master_a         (),                                                                             //    (terminated)
		.multi_ci_master_b         (),                                                                             //    (terminated)
		.multi_ci_master_c         ()                                                                              //    (terminated)
	);

	main_nios2_processor_custom_instruction_master_comb_xconnect nios2_processor_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (nios2_processor_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (nios2_processor_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (nios2_processor_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (nios2_processor_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (nios2_processor_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (nios2_processor_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (nios2_processor_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (nios2_processor_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (nios2_processor_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (nios2_processor_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (nios2_processor_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (nios2_processor_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (8),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (0)
	) nios2_processor_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (nios2_processor_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (nios2_processor_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (nios2_processor_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (nios2_processor_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (),                                                                                  // (terminated)
		.ci_master_readra    (),                                                                                  // (terminated)
		.ci_master_readrb    (),                                                                                  // (terminated)
		.ci_master_writerc   (),                                                                                  // (terminated)
		.ci_master_a         (),                                                                                  // (terminated)
		.ci_master_b         (),                                                                                  // (terminated)
		.ci_master_c         (),                                                                                  // (terminated)
		.ci_master_ipending  (),                                                                                  // (terminated)
		.ci_master_estatus   (),                                                                                  // (terminated)
		.ci_master_clk       (),                                                                                  // (terminated)
		.ci_master_clken     (),                                                                                  // (terminated)
		.ci_master_reset_req (),                                                                                  // (terminated)
		.ci_master_reset     (),                                                                                  // (terminated)
		.ci_master_start     (),                                                                                  // (terminated)
		.ci_master_done      (1'b0),                                                                              // (terminated)
		.ci_slave_clk        (1'b0),                                                                              // (terminated)
		.ci_slave_clken      (1'b0),                                                                              // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                              // (terminated)
		.ci_slave_reset      (1'b0),                                                                              // (terminated)
		.ci_slave_start      (1'b0),                                                                              // (terminated)
		.ci_slave_done       ()                                                                                   // (terminated)
	);

	main_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                       (clk_clk),                                                         //                                     clk_0_clk.clk
		.nios2_processor_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                  // nios2_processor_reset_n_reset_bridge_in_reset.reset
		.nios2_processor_data_master_address                 (nios2_processor_data_master_address),                             //                   nios2_processor_data_master.address
		.nios2_processor_data_master_waitrequest             (nios2_processor_data_master_waitrequest),                         //                                              .waitrequest
		.nios2_processor_data_master_byteenable              (nios2_processor_data_master_byteenable),                          //                                              .byteenable
		.nios2_processor_data_master_read                    (nios2_processor_data_master_read),                                //                                              .read
		.nios2_processor_data_master_readdata                (nios2_processor_data_master_readdata),                            //                                              .readdata
		.nios2_processor_data_master_write                   (nios2_processor_data_master_write),                               //                                              .write
		.nios2_processor_data_master_writedata               (nios2_processor_data_master_writedata),                           //                                              .writedata
		.nios2_processor_data_master_debugaccess             (nios2_processor_data_master_debugaccess),                         //                                              .debugaccess
		.nios2_processor_instruction_master_address          (nios2_processor_instruction_master_address),                      //            nios2_processor_instruction_master.address
		.nios2_processor_instruction_master_waitrequest      (nios2_processor_instruction_master_waitrequest),                  //                                              .waitrequest
		.nios2_processor_instruction_master_read             (nios2_processor_instruction_master_read),                         //                                              .read
		.nios2_processor_instruction_master_readdata         (nios2_processor_instruction_master_readdata),                     //                                              .readdata
		.button_down_s1_address                              (mm_interconnect_0_button_down_s1_address),                        //                                button_down_s1.address
		.button_down_s1_readdata                             (mm_interconnect_0_button_down_s1_readdata),                       //                                              .readdata
		.button_enter_s1_address                             (mm_interconnect_0_button_enter_s1_address),                       //                               button_enter_s1.address
		.button_enter_s1_write                               (mm_interconnect_0_button_enter_s1_write),                         //                                              .write
		.button_enter_s1_readdata                            (mm_interconnect_0_button_enter_s1_readdata),                      //                                              .readdata
		.button_enter_s1_writedata                           (mm_interconnect_0_button_enter_s1_writedata),                     //                                              .writedata
		.button_enter_s1_chipselect                          (mm_interconnect_0_button_enter_s1_chipselect),                    //                                              .chipselect
		.button_exit_s1_address                              (mm_interconnect_0_button_exit_s1_address),                        //                                button_exit_s1.address
		.button_exit_s1_readdata                             (mm_interconnect_0_button_exit_s1_readdata),                       //                                              .readdata
		.button_up_s1_address                                (mm_interconnect_0_button_up_s1_address),                          //                                  button_up_s1.address
		.button_up_s1_readdata                               (mm_interconnect_0_button_up_s1_readdata),                         //                                              .readdata
		.jtag_uart_0_avalon_jtag_slave_address               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),         //                 jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),           //                                              .write
		.jtag_uart_0_avalon_jtag_slave_read                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),            //                                              .read
		.jtag_uart_0_avalon_jtag_slave_readdata              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),        //                                              .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),       //                                              .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),     //                                              .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),      //                                              .chipselect
		.lcd_output_control_slave_address                    (mm_interconnect_0_lcd_output_control_slave_address),              //                      lcd_output_control_slave.address
		.lcd_output_control_slave_write                      (mm_interconnect_0_lcd_output_control_slave_write),                //                                              .write
		.lcd_output_control_slave_read                       (mm_interconnect_0_lcd_output_control_slave_read),                 //                                              .read
		.lcd_output_control_slave_readdata                   (mm_interconnect_0_lcd_output_control_slave_readdata),             //                                              .readdata
		.lcd_output_control_slave_writedata                  (mm_interconnect_0_lcd_output_control_slave_writedata),            //                                              .writedata
		.lcd_output_control_slave_begintransfer              (mm_interconnect_0_lcd_output_control_slave_begintransfer),        //                                              .begintransfer
		.led_b_s1_address                                    (mm_interconnect_0_led_b_s1_address),                              //                                      led_b_s1.address
		.led_b_s1_write                                      (mm_interconnect_0_led_b_s1_write),                                //                                              .write
		.led_b_s1_readdata                                   (mm_interconnect_0_led_b_s1_readdata),                             //                                              .readdata
		.led_b_s1_writedata                                  (mm_interconnect_0_led_b_s1_writedata),                            //                                              .writedata
		.led_b_s1_chipselect                                 (mm_interconnect_0_led_b_s1_chipselect),                           //                                              .chipselect
		.led_g_s1_address                                    (mm_interconnect_0_led_g_s1_address),                              //                                      led_g_s1.address
		.led_g_s1_write                                      (mm_interconnect_0_led_g_s1_write),                                //                                              .write
		.led_g_s1_readdata                                   (mm_interconnect_0_led_g_s1_readdata),                             //                                              .readdata
		.led_g_s1_writedata                                  (mm_interconnect_0_led_g_s1_writedata),                            //                                              .writedata
		.led_g_s1_chipselect                                 (mm_interconnect_0_led_g_s1_chipselect),                           //                                              .chipselect
		.led_r_s1_address                                    (mm_interconnect_0_led_r_s1_address),                              //                                      led_r_s1.address
		.led_r_s1_write                                      (mm_interconnect_0_led_r_s1_write),                                //                                              .write
		.led_r_s1_readdata                                   (mm_interconnect_0_led_r_s1_readdata),                             //                                              .readdata
		.led_r_s1_writedata                                  (mm_interconnect_0_led_r_s1_writedata),                            //                                              .writedata
		.led_r_s1_chipselect                                 (mm_interconnect_0_led_r_s1_chipselect),                           //                                              .chipselect
		.nios2_processor_jtag_debug_module_address           (mm_interconnect_0_nios2_processor_jtag_debug_module_address),     //             nios2_processor_jtag_debug_module.address
		.nios2_processor_jtag_debug_module_write             (mm_interconnect_0_nios2_processor_jtag_debug_module_write),       //                                              .write
		.nios2_processor_jtag_debug_module_read              (mm_interconnect_0_nios2_processor_jtag_debug_module_read),        //                                              .read
		.nios2_processor_jtag_debug_module_readdata          (mm_interconnect_0_nios2_processor_jtag_debug_module_readdata),    //                                              .readdata
		.nios2_processor_jtag_debug_module_writedata         (mm_interconnect_0_nios2_processor_jtag_debug_module_writedata),   //                                              .writedata
		.nios2_processor_jtag_debug_module_byteenable        (mm_interconnect_0_nios2_processor_jtag_debug_module_byteenable),  //                                              .byteenable
		.nios2_processor_jtag_debug_module_waitrequest       (mm_interconnect_0_nios2_processor_jtag_debug_module_waitrequest), //                                              .waitrequest
		.nios2_processor_jtag_debug_module_debugaccess       (mm_interconnect_0_nios2_processor_jtag_debug_module_debugaccess), //                                              .debugaccess
		.onchip_memory2_0_s1_address                         (mm_interconnect_0_onchip_memory2_0_s1_address),                   //                           onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                           (mm_interconnect_0_onchip_memory2_0_s1_write),                     //                                              .write
		.onchip_memory2_0_s1_readdata                        (mm_interconnect_0_onchip_memory2_0_s1_readdata),                  //                                              .readdata
		.onchip_memory2_0_s1_writedata                       (mm_interconnect_0_onchip_memory2_0_s1_writedata),                 //                                              .writedata
		.onchip_memory2_0_s1_byteenable                      (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                //                                              .byteenable
		.onchip_memory2_0_s1_chipselect                      (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                //                                              .chipselect
		.onchip_memory2_0_s1_clken                           (mm_interconnect_0_onchip_memory2_0_s1_clken),                     //                                              .clken
		.uart_main_s1_address                                (mm_interconnect_0_uart_main_s1_address),                          //                                  uart_main_s1.address
		.uart_main_s1_write                                  (mm_interconnect_0_uart_main_s1_write),                            //                                              .write
		.uart_main_s1_read                                   (mm_interconnect_0_uart_main_s1_read),                             //                                              .read
		.uart_main_s1_readdata                               (mm_interconnect_0_uart_main_s1_readdata),                         //                                              .readdata
		.uart_main_s1_writedata                              (mm_interconnect_0_uart_main_s1_writedata),                        //                                              .writedata
		.uart_main_s1_begintransfer                          (mm_interconnect_0_uart_main_s1_begintransfer),                    //                                              .begintransfer
		.uart_main_s1_chipselect                             (mm_interconnect_0_uart_main_s1_chipselect)                        //                                              .chipselect
	);

	main_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_processor_d_irq_irq)       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_processor_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (nios2_processor_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),                // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),            //          .reset_req
		.reset_req_in0  (1'b0),                                          // (terminated)
		.reset_req_in1  (1'b0),                                          // (terminated)
		.reset_in2      (1'b0),                                          // (terminated)
		.reset_req_in2  (1'b0),                                          // (terminated)
		.reset_in3      (1'b0),                                          // (terminated)
		.reset_req_in3  (1'b0),                                          // (terminated)
		.reset_in4      (1'b0),                                          // (terminated)
		.reset_req_in4  (1'b0),                                          // (terminated)
		.reset_in5      (1'b0),                                          // (terminated)
		.reset_req_in5  (1'b0),                                          // (terminated)
		.reset_in6      (1'b0),                                          // (terminated)
		.reset_req_in6  (1'b0),                                          // (terminated)
		.reset_in7      (1'b0),                                          // (terminated)
		.reset_req_in7  (1'b0),                                          // (terminated)
		.reset_in8      (1'b0),                                          // (terminated)
		.reset_req_in8  (1'b0),                                          // (terminated)
		.reset_in9      (1'b0),                                          // (terminated)
		.reset_req_in9  (1'b0),                                          // (terminated)
		.reset_in10     (1'b0),                                          // (terminated)
		.reset_req_in10 (1'b0),                                          // (terminated)
		.reset_in11     (1'b0),                                          // (terminated)
		.reset_req_in11 (1'b0),                                          // (terminated)
		.reset_in12     (1'b0),                                          // (terminated)
		.reset_req_in12 (1'b0),                                          // (terminated)
		.reset_in13     (1'b0),                                          // (terminated)
		.reset_req_in13 (1'b0),                                          // (terminated)
		.reset_in14     (1'b0),                                          // (terminated)
		.reset_req_in14 (1'b0),                                          // (terminated)
		.reset_in15     (1'b0),                                          // (terminated)
		.reset_req_in15 (1'b0)                                           // (terminated)
	);

endmodule
